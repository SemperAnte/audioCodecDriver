// full LUT tables for atan and coefd
// Automatically generated with Matlab, dont edit
localparam logic [ 63 : 0 ] atanLUTfull [ 64 ] = '{
      64'd2305843009213693952,
      64'd1361218612134873344,
      64'd719230530580880896,
      64'd365092647525521984,
      64'd183254791493294848,
      64'd91716730292036224,
      64'd45869556482713136,
      64'd22936177926750892,
      64'd11468263948075832,
      64'd5734153847876408,
      64'd2867079658191484,
      64'd1433540170878135,
      64'd716770128161890,
      64'd358385069421298,
      64'd179192535378193,
      64'd89596267772540,
      64'd44798133896700,
      64'd22399066949654,
      64'd11199533474990,
      64'd5599766737515,
      64'd2799883368760,
      64'd1399941684380,
      64'd699970842190,
      64'd349985421095,
      64'd174992710548,
      64'd87496355274,
      64'd43748177637,
      64'd21874088818,
      64'd10937044409,
      64'd5468522205,
      64'd2734261102,
      64'd1367130551,
      64'd683565276,
      64'd341782638,
      64'd170891319,
      64'd85445659,
      64'd42722830,
      64'd21361415,
      64'd10680707,
      64'd5340354,
      64'd2670177,
      64'd1335088,
      64'd667544,
      64'd333772,
      64'd166886,
      64'd83443,
      64'd41722,
      64'd20861,
      64'd10430,
      64'd5215,
      64'd2608,
      64'd1304,
      64'd652,
      64'd326,
      64'd163,
      64'd81,
      64'd41,
      64'd20,
      64'd10,
      64'd5,
      64'd3,
      64'd1,
      64'd1,
      64'd0 };

localparam logic [ 63 : 0 ] coefdLUTfull [ 26 ] = '{
      64'd3260954456333195264,
      64'd2916686334356757504,
      64'd2829601372552588288,
      64'd2807750841902562304,
      64'd2802282967498353152,
      64'd2800915666627739136,
      64'd2800573820569637376,
      64'd2800488357751430656,
      64'd2800466991965381120,
      64'd2800461650513774592,
      64'd2800460315150554624,
      64'd2800459981309729792,
      64'd2800459897849522176,
      64'd2800459876984470016,
      64'd2800459871768206848,
      64'd2800459870464141312,
      64'd2800459870138124800,
      64'd2800459870056620544,
      64'd2800459870036244480,
      64'd2800459870031150592,
      64'd2800459870029877248,
      64'd2800459870029558784,
      64'd2800459870029479424,
      64'd2800459870029459456,
      64'd2800459870029454336,
      64'd2800459870029453312 };